// This is the top level Verilog wrapper that instantiates
// the mvau.sv module. Verilog wrapper is needed for IP generation

`timescale 1ns/1ns
// Package file for parameters
 
module mvu_top #(
    parameter   KDim=2, // Kernel dimensions
    parameter   IFMCh=4,// Input feature map channels
    parameter   OFMCh=4,// Output feature map channels or the number of filter banks
    // parameter   IFMDim=4, // Input feature map dimensions
    // parameter   OFMDim=4,    // Output feature map dimensions
    parameter   SIMD=2, // Number of input columns computed in parallel
    parameter   PE=2, // Number of output rows computed in parallel
    // parameter   MMV=1, // Number of output pixels computed in parallel
    parameter   TSrcI=8, // DataType of the input activation (as used in the MAC)
    parameter   TW=1, // Word length of individual weights
    parameter   TDstI=16, // DataType of the output activation (as generated by the activation) 
    parameter   OP_SGN=0 // Enumerated values showing signedness/unsignedness of input activation/weights
//    parameter integer DSP_TRUE=0, // Use DSP blocks or LUTs for MAC
//    parameter integer INST_WMEM=1, // Instantiate weight memory, if needed
//    parameter integer MVAU_STREAM=0, // Top module is not MVAU Stream
//    parameter integer USE_ACT=0)     // Use activation after matrix-vector activation
) (    
    input           aresetn, // active low synchronous reset
    input           aclk, // main clock
    // Axis Stream interface
    input [TI-1:0]  s0_axis_tdata, // input stream
    input           s0_axis_tvalid, // input valid
    output          s0_axis_tready, // input ready
    output          m0_axis_tvalid, // output valid
    output [TO-1:0] m0_axis_tdata); // output stream
    input           m0_axis_tready, // output ready
 
mvau #(
    .KDim    (KDim      ), 
    .IFMCh   (IFMCh     ), 
    .OFMCh   (OFMCh     ), 
    .IFMDim  (IFMDim    ), 
    // .OFMDim  (OFMDim    ), 
    .SIMD    (SIMD      ), 
    .PE      (PE        ), 
    .MMV     (MMV       ), 
    .TSrcI   (TSrcI     ), 
    .TW      (TW        ), 
    .TDstI   (TDstI     ), 
    .OP_SGN  (OP_SGN    ))
mvau_inst(
    .resetn(aresetn),
    .clock(aclk),
    .rready(m0_axis_tready),
    .wready(s0_axis_tready),
    .in(s0_axis_tdata),
    .in_v(s0_axis_tvalid),
    .out_v(m0_axis_tvalid),
    .out(m0_axis_tdata)
    );
      
endmodule // mvu_top
