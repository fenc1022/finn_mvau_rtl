/*
// RTL implementation of the matrix-vector activation uint
// currently activation is not included
*/

`timescale 1ns/1ns
`include "mvu_defn.sv" // compile the package file
import mvu_defn::*; // import package into $unit compilation space

module mvu #(
    parameter int KDim=mvu_defn::KDim, // Kernel dimensions
    parameter int IFMCh=mvu_defn::IFMCh,// Input feature map channels
    parameter int OFMCh=mvu_defn::OFMCh,// Output feature map channels or the number of filter banks
    parameter int SIMD=mvu_defn::SIMD, // Number of input columns computed in parallel
    parameter int PE=mvu_defn::PE, // Number of output rows computed in parallel
    // parameter int MMV=1, // Number of output pixels computed in parallel
    parameter int TSrcI=mvu_defn::TSrcI, // DataType of the input activation (as used in the MAC)
    parameter int TW=mvu_defn::TW, // Word length of individual weights
    parameter int TDstI=mvu_defn::TDstI, // DataType of the output activation (as generated by the activation) 
    parameter bit [1:0] OP_SGN=mvu_defn::OP_SGN, // Enumerated values showing signedness/unsignedness of input activation/weights

    parameter int MatrixW=KDim*KDim*IFMCh, // Width of the input matrix
    parameter int MatrixH=OFMCh, // Heigth of the input matrix
    parameter int WMEM_DEPTH=(KDim*KDim*IFMCh*OFMCh)/(SIMD*PE), // Depth of each weight memory
    parameter int TI=SIMD*TSrcI, // SIMD times the word length of input stream
    parameter int TO=PE*TDstI // PE times the word length of output stream   
    // parameter int TA=16, // PE times the word length of the activation class (e.g thresholds)
    // parameter int DSP_TRUE=0, // Use DSP blocks or LUTs for MAC
    // parameter int INST_WMEM=1, // Instantiate weight memory, if needed
    // parameter int MVAU_STREAM=0, // Top module is not MVAU Stream
    // parameter int USE_ACT=0    // Use activation after matrix-vector activation	      
) (
    input logic             resetn,
    input logic             clock,
    // input stream
    input logic [TI-1:0]    in,
    input logic             in_v,
    output logic            wready,
    // output stream
    output logic [TO-1:0]   out,
    output logic            out_v,
    input logic             rready
);

localparam int WMEM_ADDR_BW = $clog2(WMEM_DEPTH)>1 ? $clog2(WMEM_DEPTH) : 1;
localparam int SF = MatrixW / SIMD;
localparam int NF = MatrixH / PE;

logic                    in_v_reg;
logic [TI-1:0]           in_reg;
logic [0:SIMD*TW-1]      wmem_out [0:PE-1];
logic [0:PE*SIMD*TW-1]   wmem_out_packed;
logic [TO-1:0]           out_stream;
logic                    out_stream_valid;
logic [WMEM_ADDR_BW-1:0] wmem_addr;
logic                    wmem_wready;
logic                    wmem_valid;

assign  in_v_reg = in_v;
assign  in_reg = in;

mvu_control_block #(
    .SF(SF),
    .NF(NF),
    .WMEM_DEPTH(WMEM_DEPTH))
mvu_control_block (
    .resetn,
    .clock,
    .wmem_wready,
    .wmem_valid,
    .wmem_addr
);

mvu_stream #(
    .KDim    (KDim   ),
    .IFMCh   (IFMCh  ),
    .OFMCh   (OFMCh  ),
    .MatrixW (MatrixW),
    .MatrixH (MatrixH),
    .SIMD    (SIMD   ),
    .PE      (PE     ),
    .TSrcI   (TSrcI  ),
    .TW      (TW     ),
    .TDstI   (TDstI  ),
    .OP_SGN  (OP_SGN ))
mvu_stream (
    .resetn,
    .clock,
    .in_wgt_v(wmem_valid),
    .wmem_wready,
    .in_wgt(wmem_out_packed),
    .wready,
    .in_v(in_v_reg),
    .in_act(in_reg),
    .out_v(out_stream_valid),
    .rready,
    .out(out_stream)
);

mvu_weight_mem_merged #(
    .SIMD(SIMD),
    .PE(PE),
    .TW(TW),
    .WMEM_DEPTH(WMEM_DEPTH))
mvau_weigt_mem_inst(
    .clock,
    .wmem_addr,
    .wmem_out(wmem_out)
);

generate
    for (genvar p=0; p<PE; p++)
        assign wmem_out_packed[SIMD*TW*p:SIMD*TW*(p+1)-1] = wmem_out[p];
endgenerate

logic           out_stream_valid_hold;
logic [TO-1:0]  out_stream_hold;

// Saving the 2nd stream valid if it comes
// before previous output consumed by the slave interface
always_ff @(posedge clock)
    if (!resetn)
        out_stream_valid_hold <= 1'b0;
    else if (~out_v & out_stream_valid_hold) // finish hold
        out_stream_valid_hold <= 1'b0;
    else if (out_stream_valid & out_v & ~rready)
        out_stream_valid_hold <= 1'b1;

// Saving the 2nd stream ouput if it comes
// before previous output consumed by the slave interface
always_ff @(posedge clock)
    if(!resetn)
        out_stream_hold <= 'd0;
    else if(out_stream_valid & out_v & ~rready) // Start hold
        out_stream_hold <= out_stream;

// Registered output
always_ff @(posedge clock)
    if(!resetn)
        out <= 'd0;
    else if(out_v & ~rready)
        // Hold output when input ready not asserted
        out <= out;	
    else if(out_stream_valid)
        // Read in stream unit output
        out <= out_stream; 
    else if(out_stream_valid_hold)
        // Read in the saved stream unit output which was held
        out <= out_stream_hold; 

// Output valid
always_ff @(posedge clock)
    if(!resetn) 
        out_v <= 1'b0;	    	    
    else if(out_stream_valid)
        out_v <= 1'b1;  // an output asserted by the stream unit
    else if(out_v & rready)
        out_v <= 1'b0; // output is consumed
    else if(out_stream_valid_hold)
         out_v <= 1'b1; // an output held due to non-consumption
      
endmodule