`ifndef MVAU_DEFN_PKG // if the already-compiled flag is not set
 `define MVAU_DEFN_PKG //set the flag
package mvau_defn;
   parameter VERSION = "0.1";
   parameter int KDim=2; // Kernel dimensions
   parameter int IFMCh=4;// Input feature map channels
   parameter int OFMCh=2;// Output feature map channels or the number of filter banks
   parameter int IFMDim=3; // Input feature map dimensions
   parameter int PAD=0;    // Padding around the input feature map
   parameter int STRIDE=1; // Number of pixels to move across when applying the filter
   parameter int SIMD=2; // Number of input columns computed in parallel, here SIMD < MatrixW=KDim*KDim*IFMCh
   parameter int PE=2; // Number of output rows computed in parallel, here PE <= MatrixH=OFMCh
//    parameter int WMEM_DEPTH=(KDim*KDim*IFMCh*OFMCh)/(SIMD*PE); // Depth of each weight memory
   parameter int MMV=1; // Number of output pixels computed in parallel
   parameter int TSrcI=1; // DataType of the input activation (as used in the MAC)
//    parameter int TSrcI_BIN = 0; // Indicates whether the 1-bit TSrcI is to be interpreted as special +1/-1 or not
//    parameter int TI=SIMD*TSrcI; // SIMD times the word length of input stream
   parameter int TW=1; // Word length of individual weights
//    parameter int TW_BIN = 1; // Indicates whether the 1-bit TW is to be interpreted as special +1/-1 or not
   parameter int TDstI=16; // DataType of the output activation (as generated by the activation) 
//    parameter int TA=16; // PE times the word length of the activation class (e.g thresholds)
   parameter bit [1:0] OP_SGN=2'b00; // Enumerated values showing signedness/unsignedness of input activation/weights
//    parameter int DSP_TRUE=0; // Use DSP blocks or LUTs for MAC
//    parameter int INST_WMEM=1; // Instantiate weight memory; if needed
//    parameter int USE_ACT=0;     // Use activation after matrix-vector activation
   
endpackage
   
   import mvau_defn::*; // import package into $unit compilation space
`endif
